`timescale 1ns / 1ps

//Registers 8 (Destination) contains data: 8
//Registers 20 (Source1) contains data: 10
//Registers 21 (Soruce2) contains data: 15
module PC_IM_RF(
    );

	Program_Counter PC ();
	Instruction_Memory IM ();
	Register_File ();
	

endmodule
